-- Lab 1 - ULA (S11)
-- Students: Francisco Miamoto
--           João Pedro Zanlorensi Cardoso
--           Luan Roberto
library IEEE;
use IEEE.std_logic_1164.all;

entity ula_tb is
end entity;